hi all

09-07-2023
06:22 PM
Mandya
By, Mahadevaswamy


